module cluster_level_shifter_inout (
  input  logic data_i,
  output logic data_o
);
   
  assign data_o = data_i;
   
endmodule
